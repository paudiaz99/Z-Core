
`timescale 1ns / 1ps

module axil_uart #
(
    parameter DATA_WIDTH = 32,
    parameter ADDR_WIDTH = 32,
    parameter STRB_WIDTH = (DATA_WIDTH/8)
)
(
    input  wire                   clk,
    input  wire                   rst,

    input  wire [ADDR_WIDTH-1:0]  s_axil_awaddr,
    input  wire [2:0]             s_axil_awprot,
    input  wire                   s_axil_awvalid,
    output wire                   s_axil_awready,
    input  wire [DATA_WIDTH-1:0]  s_axil_wdata,
    input  wire [STRB_WIDTH-1:0]  s_axil_wstrb,
    input  wire                   s_axil_wvalid,
    output wire                   s_axil_wready,
    output wire [1:0]             s_axil_bresp,
    output wire                   s_axil_bvalid,
    input  wire                   s_axil_bready,
    input  wire [ADDR_WIDTH-1:0]  s_axil_araddr,
    input  wire [2:0]             s_axil_arprot,
    input  wire                   s_axil_arvalid,
    output wire                   s_axil_arready,
    output wire [DATA_WIDTH-1:0]  s_axil_rdata,
    output wire [1:0]             s_axil_rresp,
    output wire                   s_axil_rvalid,
    input  wire                   s_axil_rready
);

    wire [ADDR_WIDTH-1:0] usr_addr;
    wire [DATA_WIDTH-1:0] usr_wdata;
    wire [STRB_WIDTH-1:0] usr_wstrb;
    wire usr_wen;
    wire usr_ren;
    wire [DATA_WIDTH-1:0] usr_rdata;

    assign usr_rdata = 32'h0;

    axil_slave #(
        .DATA_WIDTH(DATA_WIDTH),
        .ADDR_WIDTH(ADDR_WIDTH),
        .STRB_WIDTH(STRB_WIDTH)
    ) u_axil_slave (
        .clk(clk),
        .rst(rst),
        .s_axil_awaddr(s_axil_awaddr),
        .s_axil_awprot(s_axil_awprot),
        .s_axil_awvalid(s_axil_awvalid),
        .s_axil_awready(s_axil_awready),
        .s_axil_wdata(s_axil_wdata),
        .s_axil_wstrb(s_axil_wstrb),
        .s_axil_wvalid(s_axil_wvalid),
        .s_axil_wready(s_axil_wready),
        .s_axil_bresp(s_axil_bresp),
        .s_axil_bvalid(s_axil_bvalid),
        .s_axil_bready(s_axil_bready),
        .s_axil_araddr(s_axil_araddr),
        .s_axil_arprot(s_axil_arprot),
        .s_axil_arvalid(s_axil_arvalid),
        .s_axil_arready(s_axil_arready),
        .s_axil_rdata(s_axil_rdata),
        .s_axil_rresp(s_axil_rresp),
        .s_axil_rvalid(s_axil_rvalid),
        .s_axil_rready(s_axil_rready),
        
        // User Interface
        .usr_addr(usr_addr),
        .usr_wdata(usr_wdata),
        .usr_wstrb(usr_wstrb),
        .usr_wen(usr_wen),
        .usr_ren(usr_ren),
        .usr_rdata(usr_rdata)
    );

    // Dummy Logic for UART
    // Just acknowledge writes (handled by slave) and return 0 for reads
    // assign usr_rdata = 32'h0; // Already assigned above

    // Example: If we wanted to implement a register
    // reg [31:0] control_reg;
    // always @(posedge clk) begin
    //     if (rst) control_reg <= 0;
    //     else if (usr_wen && usr_addr[3:0] == 4'h0) control_reg <= usr_wdata;
    // end

endmodule
