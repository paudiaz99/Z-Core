module top_model (

);




endmodule