// **************************************************
//                    TODO LIST
// 1. Implement Multiple Size Load/Store
// 2. Implement AXI4 Interface
// 3. Implement Testbench (Once All Modules are Done and Tested)
// 4. Verify correctness of the Control Unit using Simulation
//
// **************************************************

`include "Core/z_core_decoder.v"
`include "Core/z_core_reg_file.v"
`include "Core/z_core_alu_ctrl.v"
`include "Core/z_core_alu.v"

module z_core_control_u 
(
    input  wire                   clk,
    input  wire                   rstn,

    output  wire [ADDR_WIDTH-1:0]  s_axil_awaddr,
    output  wire [2:0]             s_axil_awprot,
    output  wire                   s_axil_awvalid,
    input wire                   s_axil_awready,
    output wire [DATA_WIDTH-1:0]  s_axil_wdata,
    output  wire [STRB_WIDTH-1:0]  s_axil_wstrb,
    output  wire                   s_axil_wvalid,
    input wire                   s_axil_wready,
    input wire [1:0]             s_axil_bresp,
    input wire                   s_axil_bvalid,
    output wire                   s_axil_bready,
    output  wire [ADDR_WIDTH-1:0]  s_axil_araddr,
    output  wire [2:0]             s_axil_arprot,
    output  wire                   s_axil_arvalid,
    input wire                   s_axil_arready,
    input wire [DATA_WIDTH-1:0]  s_axil_rdata,
    input wire [1:0]             s_axil_rresp,
    input wire                   s_axil_rvalid,
    output wire                   s_axil_rready
);

// **************************************************
//                Instructions OP
// **************************************************

// R-Type Instructions
localparam R_INST = 7'b0110011;

// I-Type Instructions
localparam I_INST = 7'b0010011;
localparam I_LOAD_INST = 7'b0000011;
localparam JALR_INST = 7'b1100111;

// S/B-Type Instructions
localparam S_INST = 7'b0100011;
localparam B_INST = 7'b1100011;

// J/U-Type Instructions
localparam JAL_INST = 7'b1101111;
localparam LUI_INST = 7'b0110111;
localparam AUIPC_INST = 7'b0010111;

// **************************************************
//                Memory Addressing
// **************************************************

assign mem_addr = state[STATE_MEM_b] ? ALUOut_r : PC;

assign mem_write_en = state[STATE_MEM_b] ? isStore : 0;

assign mem_data_out = state[STATE_MEM_b] ? mem_data_out_r : 32'h0;

reg [31:0] MDR;
reg [31:0] mem_data_out_r;

// **************************************************
//              Instruction Register
// **************************************************

reg [31:0] IR;

// **************************************************
//                 Program Counter
// **************************************************

localparam PC_INIT = 32'd0;

// Program Counter Register
reg [31:0] PC;

// Program Counter Plus 
wire [31:0] PC_plus4     = PC + 4;
wire [31:0] PC_plus_Imm = PC + Imm_r;

// Program Counter Mux

// THIS CAN BETTER BE IMPLEMTNED USING A CASE STATEMENT
// Using a case statement, all inputs have the same propagation delay to the output
// Using nested ternary operators, the propagation delay increases with each level of nesting
// For a small number of inputs, this is not a big deal, but for a larger number of inputs, it can be significant
// Additionally, a case statement is easier to read and understand
// However, for a small number of inputs, the difference is negligible, and it comes
// down to personal preference

wire [31:0] PC_mux = (isJALR) ? alu_out :
                          isBimm           ? (alu_branch_r ? PC_plus_Imm : PC_plus4) :
                          isJAL            ? PC_plus_Imm :
                          PC_plus4;

// **************************************************
//             Instruction Decoder
// **************************************************

// Outputs
wire [6:0] op;
wire [4:0] rs1;
wire [4:0] rs2;
wire [4:0] rd;
wire [31:0] Iimm;
wire [31:0] Simm;
wire [31:0] Uimm;
wire [31:0] Bimm;
wire [31:0] Jimm;
wire [2:0] funct3;
wire [6:0] funct7;

z_core_decoder decoder (
    .inst(IR)
    ,.op(op)
    ,.rs1(rs1)
    ,.rs2(rs2)
    ,.rd(rd)
    ,.Iimm(Iimm)
    ,.Simm(Simm)
    ,.Uimm(Uimm)
    ,.Bimm(Bimm)
    ,.Jimm(Jimm)
    ,.funct3(funct3)
    ,.funct7(funct7)
);

// Decoder Combiational Logic

wire [31:0] Imm_mux_out = isIimm ? Iimm :
                          isSimm ? Simm :
                          isBimm ? Bimm :
                          isJAL  ? Jimm :
                          isUimm ? Uimm :
                          32'h0;

// Immediate Register
reg [31:0] Imm_r;

// **************************************************
//                  Register File
// **************************************************

// RD_In Multiplexer
wire [31:0] rd_in_mux = isLoad   ? MDR :
                        isJAL    ? PC_plus4 :
                        isJALR   ? PC_plus4 :
                        isLUI    ? Imm_r :
                        isAUIPC  ? PC_plus_Imm :
                        ALUOut_r;

// Outputs
wire [31:0] rs1_out;
wire [31:0] rs2_out;

z_core_reg_file reg_file (
    .clk(clk)
    ,.rd(rd)
    ,.rd_in(rd_in_mux)
    ,.rs1(rs1)
    ,.rs2(rs2)
    ,.write_enable(write_enable)
    ,.reset(~rstn)
    ,.rs1_out(rs1_out)
    ,.rs2_out(rs2_out)
);


// Write Enable Control
wire write_enable = state[STATE_WRITE_b];

// **************************************************
//                    ALU Control
// **************************************************

wire [3:0] alu_inst_type;

z_core_alu_ctrl alu_ctrl (
    .alu_op(op)
    ,.alu_funct3(funct3)
    ,.alu_funct7(funct7)
    ,.alu_inst_type(alu_inst_type)
);

// **************************************************
//                       ALU
// **************************************************

// Output Register
reg [31:0] ALUOut_r;
reg alu_branch_r;

// Outputs
wire [31:0] alu_out;
wire alu_branch;

z_core_alu alu (
    .alu_in1(alu_in1_r)
    ,.alu_in2(alu_in2_r)
    ,.alu_inst_type(alu_inst_type_r)
    ,.alu_out(alu_out)
    ,.alu_branch(alu_branch)
);

// ALU Input 2 Mux
wire [31:0] alu_in2_mux = isIimm ? Iimm :
                          isSimm ? Simm :
                          isBimm ? rs2_out :
                          isJAL  ? Jimm :
                          isUimm ? Uimm :
                          rs2_out;


// ALU Input Registers
reg [31:0] alu_in1_r;
reg [31:0] alu_in2_r;
reg [3:0] alu_inst_type_r;

// **************************************************
//                 Control Signals
// **************************************************

// Immediate Control
wire isIimm = (op == I_INST) || (op == I_LOAD_INST) || (op == JALR_INST);
wire isSimm = (op == S_INST);
wire isBimm = (op == B_INST);
wire isUimm = (op == LUI_INST) || (op == AUIPC_INST);
wire isLUI = (op == LUI_INST);
wire isAUIPC = (op == AUIPC_INST);
wire isJAL = (op == JAL_INST);
wire isJALR = (op == JALR_INST);

// Memory Control
wire isLoad = (op == I_LOAD_INST);
wire isStore = isSimm;

// WriteBack Control
wire isWB = ~(isSimm | isBimm);

// **************************************************
//                   FSM - OneHot
// **************************************************

localparam N_STATES = 5;

localparam STATE_FETCH_b   = 0;
localparam STATE_DECODE_b  = 1;
localparam STATE_EXECUTE_b = 2;
localparam STATE_MEM_b     = 3;
localparam STATE_WRITE_b   = 4;

localparam STATE_FETCH =    1 << STATE_FETCH_b;
localparam STATE_DECODE =   1 << STATE_DECODE_b;
localparam STATE_EXECUTE =  1 << STATE_EXECUTE_b;
localparam STATE_MEM =      1 << STATE_MEM_b;
localparam STATE_WRITE =    1 << STATE_WRITE_b;

reg [N_STATES-1:0] state;

always @(posedge clk) begin

    if(~rstn) begin 
        state <= STATE_FETCH;
        PC <= PC_INIT;
    end
    else begin
        if (state[STATE_FETCH_b]) begin
            // Update Instruction Register
            IR <= mem_data_in;

            state <= STATE_DECODE;
        end
        else if (state[STATE_DECODE_b]) begin
            // Update ALU Registers
            alu_in1_r <= rs1_out;
            alu_in2_r <= alu_in2_mux;
            alu_inst_type_r <= alu_inst_type;

            // Store Immediate for later use
            Imm_r <= Imm_mux_out;

            // Store rs2_out for memory store
            mem_data_out_r <= rs2_out;

            state <= STATE_EXECUTE;
        end
        else if (state[STATE_EXECUTE_b]) begin
            // Update Program Counter
            PC <= PC_mux;

            // Store ALU Results
            ALUOut_r <= alu_out;
            alu_branch_r <= alu_branch;

            state <= (isLoad || isStore) ? STATE_MEM : (isWB ? STATE_WRITE : STATE_FETCH);
        end
        else if (state[STATE_MEM_b]) begin
            // Store Memory Data Register
            if (isLoad) MDR <= mem_data_in;

            state <= isWB ? STATE_WRITE : STATE_FETCH;
        end
        else if (state[STATE_WRITE_b]) begin
            state <= STATE_FETCH;
        end
    end

end

endmodule