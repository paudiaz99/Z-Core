// **************************************************
//                    TODO LIST
// 1. Instance Control Unit, Memory, and IO Modules
// 2. Implement Testbench (Once All Modules are Done and Tested)
// 3. Verify correctness of the CPU using Simulation
// 4. Synthesize and Test on FPGA
//
// **************************************************

module top_model (

);




endmodule