// **************************************************
//                    TODO LIST
// 1. Implement Memory Controller
// 2. It has to implement a FIFO for Instruction Fetch
// 3. It has to implement a FIFO for Data Accesses
//
// **************************************************

module z_mem_controller
(
    // Inputs 

    // Outputs
);


endmodule