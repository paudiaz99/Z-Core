module z_mem_controller
(
    // Inputs 

    // Outputs
);


endmodule